-----------------------------
-- Author - Imants Pulkstenis
-- Date - 04.06.2020
-- Project name - Lab work No3
-- Module name - dds_vhdl
--
-- Detailed module description:
-- DDS sinusoidal signal generator
--
-- Revision:
-- A - initial design
-- B - 
--
-----------------------------
library ieee;					--always use this library
use ieee.std_logic_1164.all;	--always use this library

use ieee.numeric_std.all;		--use this library if arithmetic required


--define connections to outside
entity dds_vhdl is
generic
(
	phase_width 						: integer := 9;
	data_width							: integer := 16
);
port
(
	clk 								: in std_logic;	--100mhz clock
	rst									: in std_logic;	--rst
	phase_incr							: in std_Logic_vector(phase_width - 1 downto 0); --"frequency"
	phase_out							: out std_Logic_vector(phase_width - 1 downto 0);
	signal_out							: out std_Logic_vector(data_width - 1 downto 0)
);
end dds_vhdl;

--define inside of the module
architecture behavioral of dds_vhdl is

	--define inside use signals
	type rom_table is array ( 0 to 2**phase_width - 1) of std_logic_vector(data_width - 1 downto 0);
	constant signal_rom_table : rom_table := 
	(
		0 => x"0000",
		1 => x"00c9",
		2 => x"0192",
		3 => x"025b",
		4 => x"0324",
		5 => x"03ed",
		6 => x"04b5",
		7 => x"057e",
		8 => x"0646",
		9 => x"070e",
		10 => x"07d6",
		11 => x"089d",
		12 => x"0964",
		13 => x"0a2b",
		14 => x"0af1",
		15 => x"0bb7",
		16 => x"0c7c",
		17 => x"0d41",
		18 => x"0e06",
		19 => x"0eca",
		20 => x"0f8d",
		21 => x"1050",
		22 => x"1112",
		23 => x"11d3",
		24 => x"1294",
		25 => x"1354",
		26 => x"1413",
		27 => x"14d2",
		28 => x"1590",
		29 => x"164d",
		30 => x"1709",
		31 => x"17c4",
		32 => x"187e",
		33 => x"1937",
		34 => x"19f0",
		35 => x"1aa7",
		36 => x"1b5d",
		37 => x"1c12",
		38 => x"1cc7",
		39 => x"1d7a",
		40 => x"1e2b",
		41 => x"1edc",
		42 => x"1f8c",
		43 => x"203a",
		44 => x"20e7",
		45 => x"2193",
		46 => x"223e",
		47 => x"22e7",
		48 => x"238f",
		49 => x"2435",
		50 => x"24da",
		51 => x"257e",
		52 => x"2620",
		53 => x"26c1",
		54 => x"2760",
		55 => x"27fe",
		56 => x"289a",
		57 => x"2935",
		58 => x"29ce",
		59 => x"2a65",
		60 => x"2afb",
		61 => x"2b8f",
		62 => x"2c22",
		63 => x"2cb2",
		64 => x"2d41",
		65 => x"2dcf",
		66 => x"2e5a",
		67 => x"2ee4",
		68 => x"2f6c",
		69 => x"2ff2",
		70 => x"3076",
		71 => x"30f9",
		72 => x"3179",
		73 => x"31f8",
		74 => x"3274",
		75 => x"32ef",
		76 => x"3368",
		77 => x"33df",
		78 => x"3453",
		79 => x"34c6",
		80 => x"3537",
		81 => x"35a6",
		82 => x"3612",
		83 => x"367d",
		84 => x"36e5",
		85 => x"374b",
		86 => x"37b0",
		87 => x"3812",
		88 => x"3872",
		89 => x"38cf",
		90 => x"392b",
		91 => x"3984",
		92 => x"39db",
		93 => x"3a30",
		94 => x"3a83",
		95 => x"3ad3",
		96 => x"3b21",
		97 => x"3b6d",
		98 => x"3bb6",
		99 => x"3bfd",
		100 => x"3c42",
		101 => x"3c85",
		102 => x"3cc5",
		103 => x"3d03",
		104 => x"3d3f",
		105 => x"3d78",
		106 => x"3daf",
		107 => x"3de3",
		108 => x"3e15",
		109 => x"3e45",
		110 => x"3e72",
		111 => x"3e9d",
		112 => x"3ec5",
		113 => x"3eeb",
		114 => x"3f0f",
		115 => x"3f30",
		116 => x"3f4f",
		117 => x"3f6b",
		118 => x"3f85",
		119 => x"3f9c",
		120 => x"3fb1",
		121 => x"3fc4",
		122 => x"3fd4",
		123 => x"3fe1",
		124 => x"3fec",
		125 => x"3ff5",
		126 => x"3ffb",
		127 => x"3fff",
		128 => x"4000",
		129 => x"3fff",
		130 => x"3ffb",
		131 => x"3ff5",
		132 => x"3fec",
		133 => x"3fe1",
		134 => x"3fd4",
		135 => x"3fc4",
		136 => x"3fb1",
		137 => x"3f9c",
		138 => x"3f85",
		139 => x"3f6b",
		140 => x"3f4f",
		141 => x"3f30",
		142 => x"3f0f",
		143 => x"3eeb",
		144 => x"3ec5",
		145 => x"3e9d",
		146 => x"3e72",
		147 => x"3e45",
		148 => x"3e15",
		149 => x"3de3",
		150 => x"3daf",
		151 => x"3d78",
		152 => x"3d3f",
		153 => x"3d03",
		154 => x"3cc5",
		155 => x"3c85",
		156 => x"3c42",
		157 => x"3bfd",
		158 => x"3bb6",
		159 => x"3b6d",
		160 => x"3b21",
		161 => x"3ad3",
		162 => x"3a83",
		163 => x"3a30",
		164 => x"39db",
		165 => x"3984",
		166 => x"392b",
		167 => x"38cf",
		168 => x"3872",
		169 => x"3812",
		170 => x"37b0",
		171 => x"374b",
		172 => x"36e5",
		173 => x"367d",
		174 => x"3612",
		175 => x"35a6",
		176 => x"3537",
		177 => x"34c6",
		178 => x"3453",
		179 => x"33df",
		180 => x"3368",
		181 => x"32ef",
		182 => x"3274",
		183 => x"31f8",
		184 => x"3179",
		185 => x"30f9",
		186 => x"3076",
		187 => x"2ff2",
		188 => x"2f6c",
		189 => x"2ee4",
		190 => x"2e5a",
		191 => x"2dcf",
		192 => x"2d41",
		193 => x"2cb2",
		194 => x"2c22",
		195 => x"2b8f",
		196 => x"2afb",
		197 => x"2a65",
		198 => x"29ce",
		199 => x"2935",
		200 => x"289a",
		201 => x"27fe",
		202 => x"2760",
		203 => x"26c1",
		204 => x"2620",
		205 => x"257e",
		206 => x"24da",
		207 => x"2435",
		208 => x"238f",
		209 => x"22e7",
		210 => x"223e",
		211 => x"2193",
		212 => x"20e7",
		213 => x"203a",
		214 => x"1f8c",
		215 => x"1edc",
		216 => x"1e2b",
		217 => x"1d7a",
		218 => x"1cc7",
		219 => x"1c12",
		220 => x"1b5d",
		221 => x"1aa7",
		222 => x"19f0",
		223 => x"1937",
		224 => x"187e",
		225 => x"17c4",
		226 => x"1709",
		227 => x"164d",
		228 => x"1590",
		229 => x"14d2",
		230 => x"1413",
		231 => x"1354",
		232 => x"1294",
		233 => x"11d3",
		234 => x"1112",
		235 => x"1050",
		236 => x"0f8d",
		237 => x"0eca",
		238 => x"0e06",
		239 => x"0d41",
		240 => x"0c7c",
		241 => x"0bb7",
		242 => x"0af1",
		243 => x"0a2b",
		244 => x"0964",
		245 => x"089d",
		246 => x"07d6",
		247 => x"070e",
		248 => x"0646",
		249 => x"057e",
		250 => x"04b5",
		251 => x"03ed",
		252 => x"0324",
		253 => x"025b",
		254 => x"0192",
		255 => x"00c9",
		256 => x"0000",
		257 => x"ff37",
		258 => x"fe6e",
		259 => x"fda5",
		260 => x"fcdc",
		261 => x"fc13",
		262 => x"fb4b",
		263 => x"fa82",
		264 => x"f9ba",
		265 => x"f8f2",
		266 => x"f82b",
		267 => x"f763",
		268 => x"f69c",
		269 => x"f5d5",
		270 => x"f50f",
		271 => x"f449",
		272 => x"f384",
		273 => x"f2bf",
		274 => x"f1fa",
		275 => x"f136",
		276 => x"f073",
		277 => x"efb0",
		278 => x"eeee",
		279 => x"ee2d",
		280 => x"ed6c",
		281 => x"ecac",
		282 => x"ebed",
		283 => x"eb2e",
		284 => x"ea71",
		285 => x"e9b4",
		286 => x"e8f8",
		287 => x"e83c",
		288 => x"e782",
		289 => x"e6c9",
		290 => x"e611",
		291 => x"e559",
		292 => x"e4a3",
		293 => x"e3ee",
		294 => x"e33a",
		295 => x"e287",
		296 => x"e1d5",
		297 => x"e124",
		298 => x"e074",
		299 => x"dfc6",
		300 => x"df19",
		301 => x"de6d",
		302 => x"ddc3",
		303 => x"dd1a",
		304 => x"dc72",
		305 => x"dbcb",
		306 => x"db26",
		307 => x"da82",
		308 => x"d9e0",
		309 => x"d93f",
		310 => x"d8a0",
		311 => x"d802",
		312 => x"d766",
		313 => x"d6cc",
		314 => x"d633",
		315 => x"d59b",
		316 => x"d505",
		317 => x"d471",
		318 => x"d3df",
		319 => x"d34e",
		320 => x"d2bf",
		321 => x"d232",
		322 => x"d1a6",
		323 => x"d11c",
		324 => x"d094",
		325 => x"d00e",
		326 => x"cf8a",
		327 => x"cf08",
		328 => x"ce87",
		329 => x"ce09",
		330 => x"cd8c",
		331 => x"cd11",
		332 => x"cc98",
		333 => x"cc22",
		334 => x"cbad",
		335 => x"cb3a",
		336 => x"cac9",
		337 => x"ca5b",
		338 => x"c9ee",
		339 => x"c984",
		340 => x"c91b",
		341 => x"c8b5",
		342 => x"c851",
		343 => x"c7ef",
		344 => x"c78f",
		345 => x"c731",
		346 => x"c6d6",
		347 => x"c67c",
		348 => x"c625",
		349 => x"c5d0",
		350 => x"c57e",
		351 => x"c52d",
		352 => x"c4df",
		353 => x"c493",
		354 => x"c44a",
		355 => x"c403",
		356 => x"c3be",
		357 => x"c37b",
		358 => x"c33b",
		359 => x"c2fd",
		360 => x"c2c2",
		361 => x"c288",
		362 => x"c252",
		363 => x"c21d",
		364 => x"c1eb",
		365 => x"c1bb",
		366 => x"c18e",
		367 => x"c163",
		368 => x"c13b",
		369 => x"c115",
		370 => x"c0f1",
		371 => x"c0d0",
		372 => x"c0b1",
		373 => x"c095",
		374 => x"c07b",
		375 => x"c064",
		376 => x"c04f",
		377 => x"c03d",
		378 => x"c02d",
		379 => x"c01f",
		380 => x"c014",
		381 => x"c00b",
		382 => x"c005",
		383 => x"c001",
		384 => x"c000",
		385 => x"c001",
		386 => x"c005",
		387 => x"c00b",
		388 => x"c014",
		389 => x"c01f",
		390 => x"c02d",
		391 => x"c03d",
		392 => x"c04f",
		393 => x"c064",
		394 => x"c07b",
		395 => x"c095",
		396 => x"c0b1",
		397 => x"c0d0",
		398 => x"c0f1",
		399 => x"c115",
		400 => x"c13b",
		401 => x"c163",
		402 => x"c18e",
		403 => x"c1bb",
		404 => x"c1eb",
		405 => x"c21d",
		406 => x"c252",
		407 => x"c288",
		408 => x"c2c2",
		409 => x"c2fd",
		410 => x"c33b",
		411 => x"c37b",
		412 => x"c3be",
		413 => x"c403",
		414 => x"c44a",
		415 => x"c493",
		416 => x"c4df",
		417 => x"c52d",
		418 => x"c57e",
		419 => x"c5d0",
		420 => x"c625",
		421 => x"c67c",
		422 => x"c6d6",
		423 => x"c731",
		424 => x"c78f",
		425 => x"c7ef",
		426 => x"c851",
		427 => x"c8b5",
		428 => x"c91b",
		429 => x"c984",
		430 => x"c9ee",
		431 => x"ca5b",
		432 => x"cac9",
		433 => x"cb3a",
		434 => x"cbad",
		435 => x"cc22",
		436 => x"cc98",
		437 => x"cd11",
		438 => x"cd8c",
		439 => x"ce09",
		440 => x"ce87",
		441 => x"cf08",
		442 => x"cf8a",
		443 => x"d00e",
		444 => x"d094",
		445 => x"d11c",
		446 => x"d1a6",
		447 => x"d232",
		448 => x"d2bf",
		449 => x"d34e",
		450 => x"d3df",
		451 => x"d471",
		452 => x"d505",
		453 => x"d59b",
		454 => x"d633",
		455 => x"d6cc",
		456 => x"d766",
		457 => x"d802",
		458 => x"d8a0",
		459 => x"d93f",
		460 => x"d9e0",
		461 => x"da82",
		462 => x"db26",
		463 => x"dbcb",
		464 => x"dc72",
		465 => x"dd1a",
		466 => x"ddc3",
		467 => x"de6d",
		468 => x"df19",
		469 => x"dfc6",
		470 => x"e074",
		471 => x"e124",
		472 => x"e1d5",
		473 => x"e287",
		474 => x"e33a",
		475 => x"e3ee",
		476 => x"e4a3",
		477 => x"e559",
		478 => x"e611",
		479 => x"e6c9",
		480 => x"e782",
		481 => x"e83c",
		482 => x"e8f8",
		483 => x"e9b4",
		484 => x"ea71",
		485 => x"eb2e",
		486 => x"ebed",
		487 => x"ecac",
		488 => x"ed6c",
		489 => x"ee2d",
		490 => x"eeee",
		491 => x"efb0",
		492 => x"f073",
		493 => x"f136",
		494 => x"f1fa",
		495 => x"f2bf",
		496 => x"f384",
		497 => x"f449",
		498 => x"f50f",
		499 => x"f5d5",
		500 => x"f69c",
		501 => x"f763",
		502 => x"f82b",
		503 => x"f8f2",
		504 => x"f9ba",
		505 => x"fa82",
		506 => x"fb4b",
		507 => x"fc13",
		508 => x"fcdc",
		509 => x"fda5",
		510 => x"fe6e",
		511 => x"ff37"
	);
	

	-- phase counter
	signal phase_cnt : unsigned(phase_width - 1 downto 0) := (others => '0');
	



begin	--define the operation of the module!
	
	--phase output for debugging
	phase_out <= std_logic_Vector(phase_cnt);
	
	--phase counter
	process(clk)
	begin
		if rising_edge(clk) then
			if rst = '1' then		
				phase_cnt <= (others => '0');
			else
				phase_cnt <= unsigned(phase_cnt) + unsigned(phase_incr);
			end if;
		end if;
	end process;


	
	--data output
	process(clk)
	begin
		if rising_edge(clk) then
			if rst = '1' then		
				signal_out <= (others => '0');
			else
				--assign value from table
				signal_out <=  signal_rom_table(to_integer(unsigned(phase_cnt)));
			end if;
		end if;
	end process;
	
end behavioral;





